module MISO_DDR_phase_selector(
	input wire [3:0] 		phase_select,	// MISO sampling phase lag to compensate for headstage cable delay
	input wire [73:0] 	MISO4x,			// 4x oversampled MISO input
	output wire [31:0] 	MISOout				// 16-bit MISO output
	);
	
	reg[31:0] 	MISO;
	always @(*) begin
		case (phase_select)
0: MISO<={MISO4x[2],MISO4x[4],MISO4x[6],MISO4x[8],MISO4x[10],MISO4x[12],MISO4x[14],MISO4x[16],MISO4x[18],MISO4x[20],MISO4x[22],MISO4x[24],MISO4x[26],MISO4x[28],MISO4x[30],MISO4x[32],MISO4x[34],MISO4x[36],MISO4x[38],MISO4x[40],MISO4x[42],MISO4x[44],MISO4x[46],MISO4x[48],MISO4x[50],MISO4x[52],MISO4x[54],MISO4x[56],MISO4x[58],MISO4x[60],MISO4x[62]     ,MISO4x[64]};
1: MISO<={MISO4x[3],MISO4x[5],MISO4x[7],MISO4x[9],MISO4x[11],MISO4x[13],MISO4x[15],MISO4x[17],MISO4x[19],MISO4x[21],MISO4x[23],MISO4x[25],MISO4x[27],MISO4x[29],MISO4x[31],MISO4x[33],MISO4x[35],MISO4x[37],MISO4x[39],MISO4x[41],MISO4x[43],MISO4x[45],MISO4x[47],MISO4x[49],MISO4x[51],MISO4x[53],MISO4x[55],MISO4x[57],MISO4x[59],MISO4x[61],MISO4x[63]     ,MISO4x[65]};
2: MISO<={MISO4x[4],MISO4x[6],MISO4x[8],MISO4x[10],MISO4x[12],MISO4x[14],MISO4x[16],MISO4x[18],MISO4x[20],MISO4x[22],MISO4x[24],MISO4x[26],MISO4x[28],MISO4x[30],MISO4x[32],MISO4x[34],MISO4x[36],MISO4x[38],MISO4x[40],MISO4x[42],MISO4x[44],MISO4x[46],MISO4x[48],MISO4x[50],MISO4x[52],MISO4x[54],MISO4x[56],MISO4x[58],MISO4x[60],MISO4x[62],MISO4x[64]    ,MISO4x[66]};
3: MISO<={MISO4x[5],MISO4x[7],MISO4x[9],MISO4x[11],MISO4x[13],MISO4x[15],MISO4x[17],MISO4x[19],MISO4x[21],MISO4x[23],MISO4x[25],MISO4x[27],MISO4x[29],MISO4x[31],MISO4x[33],MISO4x[35],MISO4x[37],MISO4x[39],MISO4x[41],MISO4x[43],MISO4x[45],MISO4x[47],MISO4x[49],MISO4x[51],MISO4x[53],MISO4x[55],MISO4x[57],MISO4x[59],MISO4x[61],MISO4x[63],MISO4x[65]    ,MISO4x[67]};
4: MISO<={MISO4x[6],MISO4x[8],MISO4x[10],MISO4x[12],MISO4x[14],MISO4x[16],MISO4x[18],MISO4x[20],MISO4x[22],MISO4x[24],MISO4x[26],MISO4x[28],MISO4x[30],MISO4x[32],MISO4x[34],MISO4x[36],MISO4x[38],MISO4x[40],MISO4x[42],MISO4x[44],MISO4x[46],MISO4x[48],MISO4x[50],MISO4x[52],MISO4x[54],MISO4x[56],MISO4x[58],MISO4x[60],MISO4x[62],MISO4x[64],MISO4x[66]   ,MISO4x[68]};
5: MISO<={MISO4x[7],MISO4x[9],MISO4x[11],MISO4x[13],MISO4x[15],MISO4x[17],MISO4x[19],MISO4x[21],MISO4x[23],MISO4x[25],MISO4x[27],MISO4x[29],MISO4x[31],MISO4x[33],MISO4x[35],MISO4x[37],MISO4x[39],MISO4x[41],MISO4x[43],MISO4x[45],MISO4x[47],MISO4x[49],MISO4x[51],MISO4x[53],MISO4x[55],MISO4x[57],MISO4x[59],MISO4x[61],MISO4x[63],MISO4x[65],MISO4x[67]   ,MISO4x[69]};
6: MISO<={MISO4x[8],MISO4x[10],MISO4x[12],MISO4x[14],MISO4x[16],MISO4x[18],MISO4x[20],MISO4x[22],MISO4x[24],MISO4x[26],MISO4x[28],MISO4x[30],MISO4x[32],MISO4x[34],MISO4x[36],MISO4x[38],MISO4x[40],MISO4x[42],MISO4x[44],MISO4x[46],MISO4x[48],MISO4x[50],MISO4x[52],MISO4x[54],MISO4x[56],MISO4x[58],MISO4x[60],MISO4x[62],MISO4x[64],MISO4x[66],MISO4x[68]  ,MISO4x[70]};
7: MISO<={MISO4x[9],MISO4x[11],MISO4x[13],MISO4x[15],MISO4x[17],MISO4x[19],MISO4x[21],MISO4x[23],MISO4x[25],MISO4x[27],MISO4x[29],MISO4x[31],MISO4x[33],MISO4x[35],MISO4x[37],MISO4x[39],MISO4x[41],MISO4x[43],MISO4x[45],MISO4x[47],MISO4x[49],MISO4x[51],MISO4x[53],MISO4x[55],MISO4x[57],MISO4x[59],MISO4x[61],MISO4x[63],MISO4x[65],MISO4x[67],MISO4x[69]  ,MISO4x[71]};
8: MISO<={MISO4x[10],MISO4x[12],MISO4x[14],MISO4x[16],MISO4x[18],MISO4x[20],MISO4x[22],MISO4x[24],MISO4x[26],MISO4x[28],MISO4x[30],MISO4x[32],MISO4x[34],MISO4x[36],MISO4x[38],MISO4x[40],MISO4x[42],MISO4x[44],MISO4x[46],MISO4x[48],MISO4x[50],MISO4x[52],MISO4x[54],MISO4x[56],MISO4x[58],MISO4x[60],MISO4x[62],MISO4x[64],MISO4x[66],MISO4x[68],MISO4x[70] ,MISO4x[72]};
9: MISO<={MISO4x[11],MISO4x[13],MISO4x[15],MISO4x[17],MISO4x[19],MISO4x[21],MISO4x[23],MISO4x[25],MISO4x[27],MISO4x[29],MISO4x[31],MISO4x[33],MISO4x[35],MISO4x[37],MISO4x[39],MISO4x[41],MISO4x[43],MISO4x[45],MISO4x[47],MISO4x[49],MISO4x[51],MISO4x[53],MISO4x[55],MISO4x[57],MISO4x[59],MISO4x[61],MISO4x[63],MISO4x[65],MISO4x[67],MISO4x[69],MISO4x[71] ,MISO4x[73]};


default:MISO<={MISO4x[2],MISO4x[4],MISO4x[6],MISO4x[8],MISO4x[10],MISO4x[12],MISO4x[14],MISO4x[16],MISO4x[18],MISO4x[20],MISO4x[22],MISO4x[24],MISO4x[26],MISO4x[28],MISO4x[30],MISO4x[32],MISO4x[34],MISO4x[36],MISO4x[38],MISO4x[40],MISO4x[42],MISO4x[44],MISO4x[46],MISO4x[48],MISO4x[50],MISO4x[52],MISO4x[54],MISO4x[56],MISO4x[58],MISO4x[60],MISO4x[62],MISO4x[64]};
		endcase
	end

	//wire [31:0]MOSIout;
	assign MISOout[31:16]={MISO[30],MISO[28],MISO[26],MISO[24],MISO[22],MISO[20],MISO[18],MISO[16],MISO[14],MISO[12],MISO[10],MISO[8],MISO[6],MISO[4],MISO[2],MISO[0]};
	assign MISOout[15:0]={MISO[31],MISO[29],MISO[27],MISO[25],MISO[23],MISO[21],MISO[19],MISO[17],MISO[15],MISO[13],MISO[11],MISO[9],MISO[7],MISO[5],MISO[3],MISO[1]};



    endmodule